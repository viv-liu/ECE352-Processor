module FSMDecode 

endmodule
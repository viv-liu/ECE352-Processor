library verilog;
use verilog.vl_types.all;
entity multicycle_tb is
end multicycle_tb;
